
module CLK (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule

//module clock_gen(	input enable,
//						output logic clk);
//	parameter FREQ = 100000
//						
//
//endmodule : clock_gen